// Copyright (C) 2022 Intel Corporation
// SPDX-License-Identifier: MIT

`include "ofs_plat_if.vh"

//
// Top level PIM-based module.
//

module ofs_plat_afu
   (
    // All platform wires, wrapped in one interface.
    ofs_plat_if plat_ifc
    );

    // ====================================================================
    //
    //  Get an AXI-MM host channel connection from the platform.
    //
    // ====================================================================

    // Instance of the PIM's standard AXI memory interface.
    ofs_plat_axi_mem_if
      #(
        // The PIM provides parameters for configuring a standard host
        // memory DMA AXI memory interface.
        `HOST_CHAN_AXI_MEM_PARAMS,
        // PIM interfaces can be configured to log traffic during
        // simulation. In ASE, see work/log_ofs_plat_host_chan.tsv.
        .LOG_CLASS(ofs_plat_log_pkg::HOST_CHAN),

        // Set the host memory interface's burst count width so it is
        // large enough to request up to 16KB. The PIM will translate
        // large requests into sizes that are legal for the underlying
        // host channel.
        .BURST_CNT_WIDTH($clog2(16384/ofs_plat_host_chan_pkg::DATA_WIDTH_BYTES))
        )
      host_mem();

    // Instance of the PIM's AXI memory lite interface, which will be
    // used to implement the AFU's CSR space.
    ofs_plat_axi_mem_lite_if
      #(
        // The AFU choses the data bus width of the interface and the
        // PIM adjusts the address space to match.
        `HOST_CHAN_AXI_MMIO_PARAMS(64),
        // Log MMIO traffic. (See the same parameter above on host_mem.)
        .LOG_CLASS(ofs_plat_log_pkg::HOST_CHAN)
        )
        mmio64_to_afu();

    // Use the platform-provided module to map the primary host interface
    // to AXI-MM. The "primary" interface is the port that includes the
    // main OPAE-managed MMIO connection. This primary port is always
    // index 0 of plat_ifc.host_chan.ports, indepedent of the platform
    // and the native protocol of the host channel. This same module
    // name is available both on platforms that expose AXI-S PCIe TLP
    // streams to the AFU and on platforms that expose CCI-P.
    ofs_plat_host_chan_as_axi_mem_with_mmio
      #(
        // The data stream expects read responses in request order.
        // Have the PIM guarantee ordered responses. The PIM will insert
        // a reorder buffer only if read responses are not already ordered
        // by some other component, such as the PCIe SS.
        .SORT_READ_RESPONSES(1),
        // Because the algorithm in this AFU loops read responses back
        // to the host channel as writes, there is a chance for deadlocks
        // if reads and writes share ready/enable logic. No credit for
        // reads can lead to blocked writes and no way to drain pending
        // read responses. Setting BUFFER_READ_RESPONSES causes the PIM
        // to manage buffer slots for all pending read responses. If
        // the PIM has already inserted a reorder buffer the flag is
        // ignored, since the reorder buffer already has this property.
        .BUFFER_READ_RESPONSES(1)
        )
      primary_axi
       (
        .to_fiu(plat_ifc.host_chan.ports[0]),
        .host_mem_to_afu(host_mem),
        .mmio_to_afu(mmio64_to_afu),

        // These ports would be used if the PIM is told to cross to
        // a different clock. In this example, native pClk is used.
        .afu_clk(),
        .afu_reset_n()
        );


    // Each interface names its associated clock and reset.
    logic clk;
    assign clk = host_mem.clk;
    logic reset_n;
    assign reset_n = host_mem.reset_n;


    // ====================================================================
    //
    //  Get local memory from the platform.
    //
    // ====================================================================

    // The choice of interface type for local memory is independent of the
    // choice for the host channel. The host channel could be AXI-MM and
    // local memory Avalon. In fact, there is no requirement that all banks
    // of local memory be mapped to the same interface type. An AFU designer
    // who doesn't value his job could choose to map half the banks to
    // Avalon and half to AXI within a single AFU.

    ofs_plat_axi_mem_if
      #(
        `LOCAL_MEM_AXI_MEM_PARAMS_DEFAULT,
        // Log AXI transactions in simulation
        .LOG_CLASS(ofs_plat_log_pkg::LOCAL_MEM)
        )
      local_mem_to_afu[local_mem_cfg_pkg::LOCAL_MEM_NUM_BANKS]();

    // Map each bank individually
    genvar b;
    generate
        for (b = 0; b < local_mem_cfg_pkg::LOCAL_MEM_NUM_BANKS; b = b + 1)
        begin : mb
            ofs_plat_local_mem_as_axi_mem
              #(
                // Add a clock crossing from bank-specific clock.
                .ADD_CLOCK_CROSSING(1)
                )
              shim
               (
                .to_fiu(plat_ifc.local_mem.banks[b]),
                .to_afu(local_mem_to_afu[b]),

                // Map to the same clock as the AFU's host channel
                // interface. Whatever clock is chosen above in primary_hc
                // will be used here.
                .afu_clk(mmio64_to_afu.clk),
                .afu_reset_n(mmio64_to_afu.reset_n)
                );
        end
    endgenerate

    // > RP Old code TODO: Remove
    // ofs_plat_axi_mem_if
    //   #(
    //     // The PIM provides parameters for configuring a standard host
    //     // memory DMA AXI memory interface.
    //     `HOST_CHAN_AXI_MEM_PARAMS,
    //     // PIM interfaces can be configured to log traffic during
    //     // simulation. In ASE, see work/log_ofs_plat_host_chan.tsv.
    //     .LOG_CLASS(ofs_plat_log_pkg::HOST_CHAN),

    //     // Set the host memory interface's burst count width so it is
    //     // large enough to request up to 16KB. The PIM will translate
    //     // large requests into sizes that are legal for the underlying
    //     // host channel.
    //     .BURST_CNT_WIDTH($clog2(16384/ofs_plat_host_chan_pkg::DATA_WIDTH_BYTES))
    //     )
    //   ddr_mem();
    // < RP Old code TODO: Remove


    // ====================================================================
    //
    //  Tie off unused ports.
    //
    // ====================================================================

    // The PIM ties off unused devices, controlled by the AFU indicating
    // which devices it is using. This way, an AFU must know only about
    // the devices it uses. Tie-offs are thus portable, with the PIM
    // managing devices unused by and unknown to the AFU.
    ofs_plat_if_tie_off_unused
      #(
        // Host channel group 0 port 0 is connected. The mask is a
        // bit vector of indices used by the AFU.
        .HOST_CHAN_IN_USE_MASK(1),
        // All banks are used
        .LOCAL_MEM_IN_USE_MASK(-1)
        )
        tie_off(plat_ifc);


    // =========================================================================
    //
    //   Instantiate the DMA AFU.
    //
    // =========================================================================

    dma_top  
      #(
       .NUM_LOCAL_MEM_BANKS(local_mem_cfg_pkg::LOCAL_MEM_NUM_BANKS)
       )
    dma_top_inst
       (
        .mmio64_to_afu,
        .host_mem,
        .ddr_mem(local_mem_to_afu)
        );

endmodule
